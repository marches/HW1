// Simple Verilog test
module hell_test ();
initial begin
	$display("Hi");
end
endmodule